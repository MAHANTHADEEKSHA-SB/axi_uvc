class axi_transfer extends uvm_sequence_item;
   
   `uvm_object_utils(axi_transfer)
   
   function new(string name = "axi_transfer");
      super.new(name);
   endfucntion : new 
endclass : axi_transfer
