`define ADDR_WIDTH 32
`define DATA_WIDTH 32

`define ID_W_WIDTH 3
`define LOOP_W_WIDTH
`define AWCMO_WIDTH
`define BRESP_WIDTH 2

`define ID_R_WIDTH 3
`define LOOP_R_WIDTH
`define RRESP_WIDTH 2

`define USER_DATA_WIDTH
`define USER_REQ_WIDTH
`define USER_RESP_WIDTH 

`define SECSID_WIDTH
`define SID_WIDTH
`define SSID_WIDTH
`define SUBSYSID_WIDTH
`define MPAM_WIDTH
`define MECID_WIDTH 0

`define AWSNOOP_WIDTH 4
`define ARSNOOP_WIDTH 4
